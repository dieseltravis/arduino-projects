uno-music-leds
R4 3 15 220k
C2 13 0 100nF IC=0
C3 14 7 10nF IC=0
R3 12 0 10k
C1 0 15 33pF IC=0
R1 2 0 10k
C4 3 0 100nF IC=0
R2 1 0 10k

.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END
